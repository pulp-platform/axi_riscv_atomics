// Copyright (c) 2018 ETH Zurich, University of Bologna
//
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

// AXI RISC-V Atomic Operations (AMOs) Adapter
//
// This adapter implements atomic memory operations in accordance with the RVWMO memory consistency
// model.
//
// Interface notes:
// -  This module has combinational paths between AXI inputs and outputs for minimum latency. Add
//    slices upstream or downstream or in both directions if combinatorial paths become too long.
//    The module adheres to the AXI ready/valid dependency specification to prevent combinatorial
//    loops.

module axi_riscv_amos #(
    // AXI Parameters
    parameter int unsigned AXI_ADDR_WIDTH       = 0,
    parameter int unsigned AXI_DATA_WIDTH       = 0,
    parameter int unsigned AXI_ID_WIDTH         = 0,
    parameter int unsigned AXI_USER_WIDTH       = 0,
    // Maximum number of AXI write transactions outstanding at the same time
    parameter int unsigned AXI_MAX_WRITE_TXNS   = 0,
    // Word width of the widest RISC-V processor that can issue requests to this module.
    // 32 for RV32; 64 for RV64, where both 32-bit (.W suffix) and 64-bit (.D suffix) AMOs are
    // supported if `aw_strb` is set correctly.
    parameter int unsigned RISCV_WORD_WIDTH     = 0,
    /// Derived Parameters (do NOT change manually!)
    localparam int unsigned AXI_STRB_WIDTH      = AXI_DATA_WIDTH / 8
) (
    input  logic                        clk_i,
    input  logic                        rst_ni,

    /// Slave Interface
    input  logic [AXI_ADDR_WIDTH-1:0]   slv_aw_addr_i,
    input  logic [2:0]                  slv_aw_prot_i,
    input  logic [3:0]                  slv_aw_region_i,
    input  logic [5:0]                  slv_aw_atop_i,
    input  logic [7:0]                  slv_aw_len_i,
    input  logic [2:0]                  slv_aw_size_i,
    input  logic [1:0]                  slv_aw_burst_i,
    input  logic                        slv_aw_lock_i,
    input  logic [3:0]                  slv_aw_cache_i,
    input  logic [3:0]                  slv_aw_qos_i,
    input  logic [AXI_ID_WIDTH-1:0]     slv_aw_id_i,
    input  logic [AXI_USER_WIDTH-1:0]   slv_aw_user_i,
    output logic                        slv_aw_ready_o,
    input  logic                        slv_aw_valid_i,

    input  logic [AXI_ADDR_WIDTH-1:0]   slv_ar_addr_i,
    input  logic [2:0]                  slv_ar_prot_i,
    input  logic [3:0]                  slv_ar_region_i,
    input  logic [7:0]                  slv_ar_len_i,
    input  logic [2:0]                  slv_ar_size_i,
    input  logic [1:0]                  slv_ar_burst_i,
    input  logic                        slv_ar_lock_i,
    input  logic [3:0]                  slv_ar_cache_i,
    input  logic [3:0]                  slv_ar_qos_i,
    input  logic [AXI_ID_WIDTH-1:0]     slv_ar_id_i,
    input  logic [AXI_USER_WIDTH-1:0]   slv_ar_user_i,
    output logic                        slv_ar_ready_o,
    input  logic                        slv_ar_valid_i,

    input  logic [AXI_DATA_WIDTH-1:0]   slv_w_data_i,
    input  logic [AXI_STRB_WIDTH-1:0]   slv_w_strb_i,
    input  logic [AXI_USER_WIDTH-1:0]   slv_w_user_i,
    input  logic                        slv_w_last_i,
    output logic                        slv_w_ready_o,
    input  logic                        slv_w_valid_i,

    output logic [AXI_DATA_WIDTH-1:0]   slv_r_data_o,
    output logic [1:0]                  slv_r_resp_o,
    output logic                        slv_r_last_o,
    output logic [AXI_ID_WIDTH-1:0]     slv_r_id_o,
    output logic [AXI_USER_WIDTH-1:0]   slv_r_user_o,
    input  logic                        slv_r_ready_i,
    output logic                        slv_r_valid_o,

    output logic [1:0]                  slv_b_resp_o,
    output logic [AXI_ID_WIDTH-1:0]     slv_b_id_o,
    output logic [AXI_USER_WIDTH-1:0]   slv_b_user_o,
    input  logic                        slv_b_ready_i,
    output logic                        slv_b_valid_o,

    /// Master Interface
    output logic [AXI_ADDR_WIDTH-1:0]   mst_aw_addr_o,
    output logic [2:0]                  mst_aw_prot_o,
    output logic [3:0]                  mst_aw_region_o,
    output logic [5:0]                  mst_aw_atop_o,
    output logic [7:0]                  mst_aw_len_o,
    output logic [2:0]                  mst_aw_size_o,
    output logic [1:0]                  mst_aw_burst_o,
    output logic                        mst_aw_lock_o,
    output logic [3:0]                  mst_aw_cache_o,
    output logic [3:0]                  mst_aw_qos_o,
    output logic [AXI_ID_WIDTH-1:0]     mst_aw_id_o,
    output logic [AXI_USER_WIDTH-1:0]   mst_aw_user_o,
    input  logic                        mst_aw_ready_i,
    output logic                        mst_aw_valid_o,

    output logic [AXI_ADDR_WIDTH-1:0]   mst_ar_addr_o,
    output logic [2:0]                  mst_ar_prot_o,
    output logic [3:0]                  mst_ar_region_o,
    output logic [7:0]                  mst_ar_len_o,
    output logic [2:0]                  mst_ar_size_o,
    output logic [1:0]                  mst_ar_burst_o,
    output logic                        mst_ar_lock_o,
    output logic [3:0]                  mst_ar_cache_o,
    output logic [3:0]                  mst_ar_qos_o,
    output logic [AXI_ID_WIDTH-1:0]     mst_ar_id_o,
    output logic [AXI_USER_WIDTH-1:0]   mst_ar_user_o,
    input  logic                        mst_ar_ready_i,
    output logic                        mst_ar_valid_o,

    output logic [AXI_DATA_WIDTH-1:0]   mst_w_data_o,
    output logic [AXI_STRB_WIDTH-1:0]   mst_w_strb_o,
    output logic [AXI_USER_WIDTH-1:0]   mst_w_user_o,
    output logic                        mst_w_last_o,
    input  logic                        mst_w_ready_i,
    output logic                        mst_w_valid_o,

    input  logic [AXI_DATA_WIDTH-1:0]   mst_r_data_i,
    input  logic [1:0]                  mst_r_resp_i,
    input  logic                        mst_r_last_i,
    input  logic [AXI_ID_WIDTH-1:0]     mst_r_id_i,
    input  logic [AXI_USER_WIDTH-1:0]   mst_r_user_i,
    output logic                        mst_r_ready_o,
    input  logic                        mst_r_valid_i,

    input  logic [1:0]                  mst_b_resp_i,
    input  logic [AXI_ID_WIDTH-1:0]     mst_b_id_i,
    input  logic [AXI_USER_WIDTH-1:0]   mst_b_user_i,
    output logic                        mst_b_ready_o,
    input  logic                        mst_b_valid_i
);

    localparam int unsigned OUTSTND_BURSTS_WIDTH = $clog2(AXI_MAX_WRITE_TXNS+1);
    localparam int unsigned AXI_ALU_RATIO        = AXI_DATA_WIDTH/RISCV_WORD_WIDTH;

    // State types
    typedef enum logic [1:0] { FEEDTHROUGH_AW, WAIT_ALU, WAIT_AW, REQ_AW } aw_state_t;
    aw_state_t   aw_state_d, aw_state_q;

    typedef enum logic [2:0] { FEEDTHROUGH_W, WAIT_DATA, W_WAIT_RESULT, W_WAIT_CHANNEL, SEND_W } w_state_t;
    w_state_t   w_state_d, w_state_q;

    typedef enum logic [1:0] { FEEDTHROUGH_B, WAIT_B, SEND_B, VALID_REQ } b_state_t;
    b_state_t   b_state_d, b_state_q;

    typedef enum logic [1:0] { FEEDTHROUGH_AR, WAIT_AR, REQ_AR } ar_state_t;
    ar_state_t  ar_state_d, ar_state_q;

    typedef enum logic [2:0] { FEEDTHROUGH_R, WAIT_DATA_AR, CATCH_R, WAIT_R, SEND_R } r_state_t;
    r_state_t   r_state_d, r_state_q;

    typedef enum logic [1:0] { NONE, INVALID, VALID, STORE } atop_req_t;
    atop_req_t  atop_valid_d, atop_valid_q;

    // Signal declarations
    logic [OUTSTND_BURSTS_WIDTH-1:0]    w_cnt_d, w_cnt_q;
    logic [AXI_ADDR_WIDTH-1:0]          addr_d, addr_q;
    logic [AXI_ID_WIDTH-1:0]            id_d, id_q;
    logic [2:0]                         size_d, size_q;
    logic [AXI_STRB_WIDTH-1:0]          strb_d, strb_q;
    logic [3:0]                         cache_d, cache_q;
    logic [2:0]                         prot_d, prot_q;
    logic [3:0]                         qos_d, qos_q;
    logic [3:0]                         region_d, region_q;
    logic [AXI_USER_WIDTH-1:0]          user_d, user_q;
    logic [AXI_DATA_WIDTH-1:0]          atop_data_d, atop_data_q;
    logic [AXI_DATA_WIDTH-1:0]          read_data_d, read_data_q;
    logic [AXI_DATA_WIDTH-1:0]          write_data_d, write_data_q;
    logic [5:0]                         atop_d, atop_q;
    logic                               data_valid_d, data_valid_q;

    logic                               read_done_d, read_done_q;
    logic                               adapter_ready;

    logic [RISCV_WORD_WIDTH-1:0]    alu_operand_a;
    logic [RISCV_WORD_WIDTH-1:0]    alu_operand_b;
    logic [RISCV_WORD_WIDTH-1:0]    alu_result;
    logic [AXI_DATA_WIDTH-1:0]      alu_result_ext;

    /**
     * Calculate ready signals and channel states
     */

    // Check if all state machines are ready for the next atomic request
    assign adapter_ready = (aw_state_q == FEEDTHROUGH_AW) &&
                           ( w_state_q == FEEDTHROUGH_W ) &&
                           ( b_state_q == FEEDTHROUGH_B ) &&
                           (ar_state_q == FEEDTHROUGH_AR) &&
                           ( r_state_q == FEEDTHROUGH_R );

    // Calculate if the channels are free
    logic aw_valid, aw_ready;
    logic  w_valid,  w_ready;
    logic  b_valid,  b_ready;
    logic ar_valid, ar_ready;
    logic  r_valid,  r_ready;
    logic aw_free, w_free, b_free, ar_free, r_free;

    assign aw_free = ~aw_valid | aw_ready;
    assign  w_free = ~ w_valid |  w_ready;
    assign  b_free = ~ b_valid |  b_ready;
    assign ar_free = ~ar_valid | ar_ready;
    assign  r_free = ~ r_valid |  r_ready;

    always_ff @(posedge clk_i or negedge rst_ni) begin
        if(~rst_ni) begin
            aw_valid <= 0;
            aw_ready <= 0;
            w_valid  <= 0;
            w_ready  <= 0;
            b_valid  <= 0;
            b_ready  <= 0;
            ar_valid <= 0;
            ar_ready <= 0;
            r_valid  <= 0;
            r_ready  <= 0;
        end else begin
            aw_valid <= mst_aw_valid_o;
            aw_ready <= mst_aw_ready_i;
            w_valid  <= mst_w_valid_o;
            w_ready  <= mst_w_ready_i;
            b_valid  <= slv_b_valid_o;
            b_ready  <= slv_b_ready_i;
            ar_valid <= mst_ar_valid_o;
            ar_ready <= mst_ar_ready_i;
            r_valid  <= slv_r_valid_o;
            r_ready  <= slv_r_ready_i;
        end
    end

    // Calculate if the request interferes with the ongoing atomic transaction
    // The protected bytes go from addr_q up to addr_q + (1 << size_q) - 1
    // TODO Bursts need special treatment
    // TODO Some memory controller round the address down
    logic transaction_collision;
    assign transaction_collision = (slv_aw_addr_i < (     addr_q + (8'h01 <<      size_q))) &
                                   (     addr_q < (slv_aw_addr_i + (8'h01 << slv_aw_size_i)));

    always_comb begin : calc_atop_valid
        atop_valid_d = atop_valid_q;
        if (adapter_ready) begin
            atop_valid_d = NONE;
            if (slv_aw_valid_i && slv_aw_atop_i) begin
                // Default is invalid request
                atop_valid_d = INVALID;
                // Valid load operation
                if ((slv_aw_atop_i      ==  axi_pkg::ATOP_ATOMICSWAP) ||
                    (slv_aw_atop_i[5:3] == {axi_pkg::ATOP_ATOMICLOAD , axi_pkg::ATOP_LITTLE_END})) begin
                    atop_valid_d = VALID;
                end
                // Valid store operation
                if (slv_aw_atop_i[5:3] == {axi_pkg::ATOP_ATOMICSTORE, axi_pkg::ATOP_LITTLE_END}) begin
                    atop_valid_d = STORE;
                end
                // Invalidate valid request if control signals do not match
                // Burst or exclusive access
                if (slv_aw_len_i | slv_aw_lock_i) begin
                    atop_valid_d = INVALID;
                end
                // Unsupported size
                if (slv_aw_size_i > $clog2(RISCV_WORD_WIDTH/8)) begin
                    atop_valid_d = INVALID;
                end
            end
        end
    end

    always_ff @(posedge clk_i or negedge rst_ni) begin : proc_atop_valid
        if(~rst_ni) begin
            atop_valid_q <= NONE;
        end else begin
            atop_valid_q <= atop_valid_d;
        end
    end

    /**
     * Write Channel: AW, W, B
     */

    /*====================================================================
    =                                 AW                                 =
    ====================================================================*/
    logic [OUTSTND_BURSTS_WIDTH-1:0]  w_cnt_inj_d, w_cnt_inj_q;

    always_comb begin : axi_aw_channel
        // Defaults
        mst_aw_id_o     = slv_aw_id_i;
        mst_aw_addr_o   = slv_aw_addr_i;
        mst_aw_len_o    = slv_aw_len_i;
        mst_aw_size_o   = slv_aw_size_i;
        mst_aw_burst_o  = slv_aw_burst_i;
        mst_aw_lock_o   = slv_aw_lock_i;
        mst_aw_cache_o  = slv_aw_cache_i;
        mst_aw_prot_o   = slv_aw_prot_i;
        mst_aw_qos_o    = slv_aw_qos_i;
        mst_aw_region_o = slv_aw_region_i;
        mst_aw_atop_o   = 6'b0;
        mst_aw_user_o   = slv_aw_user_i;
        // Non-AXI signals
        addr_d       = addr_q;
        id_d         = id_q;
        size_d       = size_q;
        atop_d       = atop_q;
        cache_d      = cache_q;
        prot_d       = prot_q;
        qos_d        = qos_q;
        region_d     = region_q;
        user_d       = user_q;
        w_cnt_inj_d  = w_cnt_inj_q;
        // State Machine
        aw_state_d   = aw_state_q;

        // Default control
        // Make sure the outstanding beats counter does not overflow
        if (w_cnt_q == AXI_MAX_WRITE_TXNS || (slv_aw_valid_i && slv_aw_atop_i)) begin
            // Block if counter is overflowing or atomic request
            mst_aw_valid_o = 1'b0;
            slv_aw_ready_o = 1'b0;
        end else if (slv_aw_valid_i && transaction_collision && !adapter_ready) begin
            // Block requests to the same address as current atomic transaction
            mst_aw_valid_o = 1'b0;
            slv_aw_ready_o = 1'b0;
        end else begin
            // Forward
            mst_aw_valid_o  = slv_aw_valid_i;
            slv_aw_ready_o  = mst_aw_ready_i;
        end

        unique case (aw_state_q)

            FEEDTHROUGH_AW: begin
                // Feedthrough slave to master until atomic operation is detected
                if (slv_aw_valid_i && slv_aw_atop_i) begin
                    // Do not forward
                    mst_aw_valid_o = 1'b0;
                    if (adapter_ready) begin
                        // Acknowledge atomic transaction
                        slv_aw_ready_o = 1'b1;
                        // Remember request
                        atop_d   = slv_aw_atop_i;
                        addr_d   = slv_aw_addr_i;
                        id_d     = slv_aw_id_i;
                        size_d   = slv_aw_size_i;
                        cache_d  = slv_aw_cache_i;
                        prot_d   = slv_aw_prot_i;
                        qos_d    = slv_aw_qos_i;
                        region_d = slv_aw_region_i;
                        user_d   = slv_aw_user_i;
                        // Go to next state
                        if (atop_valid_d != INVALID) begin
                            aw_state_d = WAIT_ALU;
                        end
                    end else begin
                        // Block request
                        slv_aw_ready_o  = 1'b0;
                    end
                end

                // Keep counting the W beats
                if (w_cnt_inj_q && mst_w_valid_o && mst_w_ready_i && mst_w_last_o) begin
                    w_cnt_inj_d = w_cnt_inj_q - 1;
                end
            end // FEEDTHROUGH_AW

            WAIT_ALU: begin
                w_cnt_inj_d = 1'b0;
                // If the result is ready, try to write it
                if (read_done_q && data_valid_q) begin
                    // Check if AW channel is free
                    if (aw_free) begin
                        // Block
                        slv_aw_ready_o  = 1'b0;
                        // Make write request
                        mst_aw_valid_o  = 1'b1;
                        mst_aw_addr_o   = addr_q;
                        mst_aw_len_o    = 8'h00;
                        mst_aw_id_o     = id_q;
                        mst_aw_size_o   = size_q;
                        mst_aw_burst_o  = 2'b00;
                        mst_aw_lock_o   = 1'b0;
                        mst_aw_cache_o  = cache_q;
                        mst_aw_prot_o   = prot_q;
                        mst_aw_qos_o    = qos_q;
                        mst_aw_region_o = region_q;
                        mst_aw_user_o   = user_q;
                        // Remember outstanding beats before injected request
                        if (mst_w_valid_o && mst_w_ready_i && mst_w_last_o) begin
                            w_cnt_inj_d = w_cnt_q - 1;
                        end else begin
                            w_cnt_inj_d = w_cnt_q;
                        end
                        // Check if request is acknowledged
                        if (mst_aw_ready_i) begin
                            aw_state_d = FEEDTHROUGH_AW;
                        end else begin
                            aw_state_d = REQ_AW;
                        end
                    end else begin
                    end
                end
            end // WAIT_ALU

            REQ_AW: begin
                // Block
                slv_aw_ready_o  = 1'b0;
                // Hold write request
                mst_aw_valid_o  = 1'b1;
                mst_aw_addr_o   = addr_q;
                mst_aw_len_o    = 8'h00;
                mst_aw_id_o     = id_q;
                mst_aw_size_o   = size_q;
                mst_aw_burst_o  = 2'b00;
                mst_aw_lock_o   = 1'b0;
                mst_aw_cache_o  = cache_q;
                mst_aw_prot_o   = prot_q;
                mst_aw_qos_o    = qos_q;
                mst_aw_region_o = region_q;
                mst_aw_user_o   = user_q;
                if (mst_aw_ready_i) begin
                    aw_state_d = FEEDTHROUGH_AW;
                end
                // Keep counting the W beats
                if (w_cnt_inj_q && mst_w_valid_o && mst_w_ready_i && mst_w_last_o) begin
                    w_cnt_inj_d = w_cnt_inj_q - 1;
                end
            end // REQ_AW

            default: aw_state_d = FEEDTHROUGH_AW;

        endcase
    end // axi_aw_channel

    /*====================================================================
    =                                 W                                  =
    ====================================================================*/
    logic [OUTSTND_BURSTS_WIDTH-1:0]  w_cnt_req_d, w_cnt_req_q;

    always_comb begin : axi_w_channel
        // Defaults
        mst_w_data_o = slv_w_data_i;
        mst_w_strb_o = slv_w_strb_i;
        mst_w_last_o = slv_w_last_i;
        mst_w_user_o = slv_w_user_i;
        // Non-AXI signals
        strb_d       = strb_q;
        atop_data_d  = atop_data_q;
        write_data_d = write_data_q;
        data_valid_d = data_valid_q;
        // State Machine
        w_state_d   = w_state_q;
        w_cnt_req_d = w_cnt_req_q;

        // Default control
        // Make sure no data is sent without knowing if it's atomic
        if (w_cnt_q == 0) begin
            // Stall W as it precedes the AW request
            slv_w_ready_o = 1'b0;
            mst_w_valid_o = 1'b0;
        end else begin
            mst_w_valid_o = slv_w_valid_i;
            slv_w_ready_o = mst_w_ready_i;
        end

        unique case (w_state_q)

            FEEDTHROUGH_W: begin
                if (adapter_ready) begin
                    // Reset read flag
                    data_valid_d = 1'b0;
                    write_data_d = '0;

                    if (atop_valid_d != NONE) begin
                        // Check if data is also available and does not belong to previous request
                        if (w_cnt_q == 0) begin
                            // Block downstream
                            mst_w_valid_o = 1'b0;
                            // Fetch data and wait for all data
                            slv_w_ready_o  = 1'b1;
                            if (slv_w_valid_i) begin
                                if (atop_valid_d != INVALID) begin
                                    atop_data_d  = slv_w_data_i;
                                    strb_d       = slv_w_strb_i;
                                    data_valid_d = 1'b1;
                                    w_state_d    = W_WAIT_RESULT;
                                end
                            end else begin
                                w_cnt_req_d = '0;
                                w_state_d   = WAIT_DATA;
                            end
                        end else begin
                            // Remember the amount of outstanding bursts and count down
                            if (mst_w_valid_o && mst_w_ready_i && mst_w_last_o) begin
                                w_cnt_req_d = w_cnt_q - 1;
                            end else begin
                                w_cnt_req_d = w_cnt_q;
                            end
                            w_state_d   = WAIT_DATA;
                        end
                    end
                end
            end // FEEDTHROUGH_W

            WAIT_DATA: begin
                // Count W beats until data arrives that belongs to the AMO request
                if (w_cnt_req_q == 0) begin
                    // Block downstream
                    mst_w_valid_o = 1'b0;
                    // Ready upstream
                    slv_w_ready_o = 1'b1;

                    if (slv_w_valid_i) begin
                        if (atop_valid_q == INVALID) begin
                            w_state_d    = FEEDTHROUGH_W;
                        end else begin
                            atop_data_d  = slv_w_data_i;
                            strb_d       = slv_w_strb_i;
                            data_valid_d = 1'b1;
                            w_state_d    = W_WAIT_RESULT;
                        end
                    end
                end else if (mst_w_valid_o && mst_w_ready_i && mst_w_last_o) begin
                    w_cnt_req_d = w_cnt_req_q - 1;
                end
            end

            W_WAIT_RESULT: begin
                // If the result is ready, try to write it
                if (read_done_q && data_valid_q && aw_free) begin
                    // Check if W channel is free and make sure data is not interleaved
                    write_data_d = alu_result_ext;
                    if (w_free && w_cnt_q == 0) begin
                        // Block
                        slv_w_ready_o  = 1'b0;
                        // Send write data
                        mst_w_valid_o  = 1'b1;
                        mst_w_data_o   = alu_result_ext;
                        mst_w_last_o   = 1'b1;
                        mst_w_strb_o   = strb_q;
                        if (mst_w_ready_i) begin
                            w_state_d = FEEDTHROUGH_W;
                        end else begin
                            w_state_d = SEND_W;
                        end
                    end else begin
                        w_state_d = W_WAIT_CHANNEL;
                    end
                end
            end // W_WAIT_RESULT

            W_WAIT_CHANNEL: begin
                // Wait to not interleave the data
                if (w_free && w_cnt_inj_q == 0) begin
                    // Block
                    slv_w_ready_o = 1'b0;
                    // Send write data
                    mst_w_valid_o  = 1'b1;
                    mst_w_data_o   = write_data_q;
                    mst_w_last_o   = 1'b1;
                    mst_w_strb_o   = strb_q;
                    if (mst_w_ready_i) begin
                        w_state_d = FEEDTHROUGH_W;
                    end else begin
                        w_state_d = SEND_W;
                    end
                end
            end // W_WAIT_CHANNEL

            SEND_W: begin
                // Block
                slv_w_ready_o = 1'b0;
                // Send write data
                mst_w_valid_o  = 1'b1;
                mst_w_data_o   = write_data_q;
                mst_w_last_o   = 1'b1;
                mst_w_strb_o   = strb_q;
                if (mst_w_ready_i) begin
                    w_state_d = FEEDTHROUGH_W;
                end
            end // SEND_W

            default: w_state_d = FEEDTHROUGH_W;

        endcase
    end // axi_w_channel

    /*====================================================================
    =                                 B                                  =
    ====================================================================*/
    always_comb begin : axi_b_channel
        // Defaults
        mst_b_ready_o  = slv_b_ready_i;
        slv_b_id_o     = mst_b_id_i;
        slv_b_resp_o   = mst_b_resp_i;
        slv_b_user_o   = mst_b_user_i;
        slv_b_valid_o  = mst_b_valid_i;
        // State Machine
        b_state_d    = b_state_q;

        unique case (b_state_q)

            FEEDTHROUGH_B: begin
                if (adapter_ready) begin
                    if (atop_valid_d == VALID || atop_valid_d == STORE) begin
                        b_state_d = VALID_REQ;
                    end else if (atop_valid_d == INVALID) begin
                        // Inject B resp
                        // Check if the B channel is free
                        if (mst_b_valid_i) begin
                            b_state_d   = WAIT_B;
                        end else begin
                            mst_b_ready_o  = 1'b0;
                            // Write B response
                            slv_b_id_o     = slv_aw_id_i;
                            slv_b_resp_o   = axi_pkg::RESP_SLVERR;
                            slv_b_valid_o  = 1'b1;
                            if (!slv_b_ready_i) begin
                                b_state_d = SEND_B;
                            end
                        end
                    end
                end
            end // FEEDTHROUGH_B

            WAIT_B, SEND_B: begin
                if (b_free || (b_state_q == SEND_B)) begin
                    mst_b_ready_o  = 1'b0;
                    // Write B response
                    slv_b_id_o     = id_q;
                    slv_b_resp_o   = axi_pkg::RESP_SLVERR;
                    slv_b_valid_o  = 1'b1;
                    if (slv_b_ready_i) begin
                        b_state_d = FEEDTHROUGH_B;
                    end else begin
                        b_state_d = SEND_B;
                    end
                end
            end // WAIT_B

            VALID_REQ: begin
                if (mst_b_valid_i && mst_b_id_i == id_q) begin
                    b_state_d = FEEDTHROUGH_B;
                end
            end // VALID_REQ

            default: b_state_d = FEEDTHROUGH_B;

        endcase
    end // axi_b_channel

    // Keep track of outstanding downstream write bursts and responses.
    always_comb begin
        w_cnt_d = w_cnt_q;
        if (mst_aw_valid_o && mst_aw_ready_i) begin
            w_cnt_d += 1;
        end
        if (mst_w_valid_o && mst_w_ready_i && mst_w_last_o) begin
            w_cnt_d -= 1;
        end
    end

    always_ff @(posedge clk_i or negedge rst_ni) begin : axi_write_channel_ff
        if(~rst_ni) begin
            aw_state_q   <= FEEDTHROUGH_AW;
            w_state_q    <= FEEDTHROUGH_W;
            b_state_q    <= FEEDTHROUGH_B;
            w_cnt_q      <= '0;
            w_cnt_req_q  <= '0;
            w_cnt_inj_q  <= '0;
            addr_q       <= '0;
            id_q         <= '0;
            size_q       <= '0;
            strb_q       <= '0;
            cache_q      <= '0;
            prot_q       <= '0;
            qos_q        <= '0;
            region_q     <= '0;
            user_q       <= '0;
            atop_data_q  <= '0;
            write_data_q <= '0;
            data_valid_q <= '0;
            atop_q       <= 6'b0;
        end else begin
            aw_state_q   <= aw_state_d;
            w_state_q    <= w_state_d;
            b_state_q    <= b_state_d;
            w_cnt_q      <= w_cnt_d;
            w_cnt_req_q  <= w_cnt_req_d;
            w_cnt_inj_q  <= w_cnt_inj_d;
            addr_q       <= addr_d;
            id_q         <= id_d;
            size_q       <= size_d;
            strb_q       <= strb_d;
            cache_q      <= cache_d;
            prot_q       <= prot_d;
            qos_q        <= qos_d;
            region_q     <= region_d;
            user_q       <= user_d;
            atop_data_q  <= atop_data_d;
            write_data_q <= write_data_d;
            data_valid_q <= data_valid_d;
            atop_q       <= atop_d;
        end
    end

    /**
    * Read Channel: AR, R
    */

    /*====================================================================
    =                                AR                                  =
    ====================================================================*/
    always_comb begin : axi_AR_channel
        mst_ar_id_o     = slv_ar_id_i;
        mst_ar_addr_o   = slv_ar_addr_i;
        mst_ar_len_o    = slv_ar_len_i;
        mst_ar_size_o   = slv_ar_size_i;
        mst_ar_burst_o  = slv_ar_burst_i;
        mst_ar_lock_o   = slv_ar_lock_i;
        mst_ar_cache_o  = slv_ar_cache_i;
        mst_ar_prot_o   = slv_ar_prot_i;
        mst_ar_qos_o    = slv_ar_qos_i;
        mst_ar_region_o = slv_ar_region_i;
        mst_ar_user_o   = slv_ar_user_i;
        mst_ar_valid_o  = 1'b0;
        slv_ar_ready_o  = 1'b0;

        // State Machine
        ar_state_d  = ar_state_q;

        unique case (ar_state_q)

            FEEDTHROUGH_AR: begin
                // Feed through
                mst_ar_valid_o  = slv_ar_valid_i;
                slv_ar_ready_o  = mst_ar_ready_i;

                if (adapter_ready) begin
                    if (atop_valid_d == VALID | atop_valid_d == STORE) begin
                        if (slv_ar_valid_i) begin
                            // Wait until AR is free
                            ar_state_d   = WAIT_AR;
                        end else begin
                            // Acquire channel
                            slv_ar_ready_o  = 1'b0;
                            // Immediately start read request
                            mst_ar_addr_o   = slv_aw_addr_i;
                            mst_ar_id_o     = slv_aw_id_i;
                            mst_ar_len_o    = 8'h00;
                            mst_ar_size_o   = slv_aw_size_i;
                            mst_ar_burst_o  = 2'b00;
                            mst_ar_lock_o   = 1'h0;
                            mst_ar_valid_o  = 1'b1;
                            if (!mst_ar_ready_i) begin
                                // Hold read request but do not depend on AW
                                ar_state_d = REQ_AR;
                            end
                        end
                    end
                end
            end // FEEDTHROUGH_AR

            WAIT_AR: begin
                // Issue read request
                if (ar_free) begin
                    // Inject read request
                    mst_ar_addr_o   = addr_q;
                    mst_ar_id_o     = id_q;
                    mst_ar_len_o    = 8'h00;
                    mst_ar_size_o   = size_q;
                    mst_ar_burst_o  = 2'b00;
                    mst_ar_lock_o   = 1'h0;
                    mst_ar_valid_o  = 1'b1;
                    if (mst_ar_ready_i) begin
                        // Request acknowledged
                        ar_state_d = FEEDTHROUGH_AR;
                    end else begin
                        // Hold read request
                        ar_state_d = REQ_AR;
                    end
                end else begin
                    // Wait until AR is free
                    mst_ar_valid_o = slv_ar_valid_i;
                    slv_ar_ready_o = mst_ar_ready_i;
                end
            end // WAIT_AR

            REQ_AR: begin
                // Inject read request
                mst_ar_addr_o   = addr_q;
                mst_ar_id_o     = id_q;
                mst_ar_len_o    = 8'h00;
                mst_ar_size_o   = size_q;
                mst_ar_burst_o  = 2'b00;
                mst_ar_lock_o   = 1'h0;
                mst_ar_valid_o  = 1'b1;
                if (mst_ar_ready_i) begin
                    // Request acknowledged
                    ar_state_d = FEEDTHROUGH_AR;
                end
            end // REQ_AR

            default: ar_state_d = FEEDTHROUGH_AR;

        endcase
    end

    /*====================================================================
    =                                 R                                  =
    ====================================================================*/
    always_comb begin : axi_R_channel

        // Feed through the R channel by default
        mst_r_ready_o   = slv_r_ready_i;
        slv_r_id_o      = mst_r_id_i;
        slv_r_data_o    = mst_r_data_i;
        slv_r_resp_o    = mst_r_resp_i;
        slv_r_last_o    = mst_r_last_i;
        slv_r_user_o    = mst_r_user_i;
        slv_r_valid_o   = mst_r_valid_i;

        // State Machine
        read_data_d = read_data_q;
        read_done_d = read_done_q;
        r_state_d   = r_state_q;

        unique case (r_state_q)

            FEEDTHROUGH_R: begin
                if (adapter_ready) begin
                    // Reset read flag
                    read_done_d  = 1'b0;

                    if (atop_valid_d == VALID) begin
                        // Wait for R response to read data
                        r_state_d = WAIT_DATA_AR;
                    end else if (atop_valid_d == INVALID) begin
                        // Send R response
                        // Check if the R channel is free
                        if (mst_r_valid_i) begin
                            r_state_d = WAIT_R;
                        end else begin
                            // Acquire the R channel
                            slv_r_valid_o = 1'b0;
                            mst_r_ready_o = 1'b0;
                            r_state_d   = SEND_R;
                        end
                    end else if (atop_valid_d == STORE) begin
                        // Wait for R response to catch
                        r_state_d = CATCH_R;
                    end
                end
            end // FEEDTHROUGH_R

            WAIT_DATA_AR: begin
                // Read data
                if (mst_r_valid_i && (mst_r_id_i == id_q)) begin
                    read_data_d = mst_r_data_i;
                    read_done_d = 1'b1;
                    if (slv_r_ready_i) begin
                        r_state_d  = FEEDTHROUGH_R;
                    end
                end
            end // WAIT_DATA_AR

            CATCH_R: begin
                // Atomic store --> block the R response
                if (mst_r_valid_i && (mst_r_id_i == id_q)) begin
                    // Block
                    slv_r_valid_o = 1'b0;
                    // ACK
                    mst_r_ready_o = 1'b1;
                    // Store data
                    read_data_d = mst_r_data_i;
                    read_done_d = 1'b1;
                    r_state_d   = FEEDTHROUGH_R;
                end
            end // CATCH_R

            WAIT_R: begin
                // Wait for the R channel to become free
                if (r_free) begin
                    // Block memory
                    mst_r_ready_o = 1'b0;
                    // Send own R resp
                    slv_r_valid_o = 1'b1;
                    slv_r_data_o  = '1;
                    slv_r_id_o    = id_q;
                    slv_r_resp_o  = axi_pkg::RESP_SLVERR;
                    slv_r_last_o  = 1'b1;
                    if (slv_r_ready_i) begin
                        r_state_d = FEEDTHROUGH_R;
                    end else begin
                        r_state_d = SEND_R;
                    end
                end
            end // WAIT_R

            SEND_R: begin
                // Block memory
                mst_r_ready_o = 1'b0;
                // Send own R resp
                slv_r_valid_o = 1'b1;
                slv_r_data_o  = '1;
                slv_r_id_o    = id_q;
                slv_r_resp_o  = axi_pkg::RESP_SLVERR;
                slv_r_last_o  = 1'b1;
                if (slv_r_ready_i) begin
                    r_state_d = FEEDTHROUGH_R;
                end
            end // SEND_R

            default: r_state_d = FEEDTHROUGH_R;

        endcase
    end

    always_ff @(posedge clk_i or negedge rst_ni) begin : axi_read_channel_ff
        if(~rst_ni) begin
            ar_state_q  <= FEEDTHROUGH_AR;
            r_state_q   <= FEEDTHROUGH_R;
            read_data_q <= '0;
            read_done_q <= 1'b0;
        end else begin
            ar_state_q  <= ar_state_d;
            r_state_q   <= r_state_d;
            read_data_q <= read_data_d;
            read_done_q <= read_done_d;
        end
    end

    /**
     * ALU
     */

    logic [AXI_ALU_RATIO-1:0][RISCV_WORD_WIDTH-1:0] op_a;
    logic [AXI_ALU_RATIO-1:0][RISCV_WORD_WIDTH-1:0] op_b;
    logic [AXI_ALU_RATIO-1:0][RISCV_WORD_WIDTH-1:0] op_a_sign_ext;
    logic [AXI_ALU_RATIO-1:0][RISCV_WORD_WIDTH-1:0] op_b_sign_ext;
    logic [AXI_ALU_RATIO-1:0][RISCV_WORD_WIDTH-1:0] res;
    logic [AXI_STRB_WIDTH-1:0][7:0]                 strb_ext;
    logic sign_a;
    logic sign_b;

    assign op_a = read_data_q & strb_ext;
    assign op_b = atop_data_q & strb_ext;
    assign sign_a = |(op_a & ~(strb_ext >> 1));
    assign sign_b = |(op_b & ~(strb_ext >> 1));
    assign alu_result_ext = res;

    generate
        if (AXI_ALU_RATIO == 1 && RISCV_WORD_WIDTH == 32) begin
            assign alu_operand_a  = op_a;
            assign alu_operand_b  = op_b;
            assign res            = alu_result;
        end else if (AXI_ALU_RATIO == 1 && RISCV_WORD_WIDTH == 64) begin
            assign res        = alu_result;
            always_comb begin
                op_a_sign_ext = op_a | ({AXI_ALU_RATIO*RISCV_WORD_WIDTH{sign_a}} & ~strb_ext);
                op_b_sign_ext = op_b | ({AXI_ALU_RATIO*RISCV_WORD_WIDTH{sign_b}} & ~strb_ext);

                if (atop_q[2:0] == axi_pkg::ATOP_SMAX || atop_q[2:0] == axi_pkg::ATOP_SMIN) begin
                    // Sign extend
                    alu_operand_a = op_a_sign_ext;
                    alu_operand_b = op_b_sign_ext;
                end else begin
                    // No sign extension necessary
                    alu_operand_a = op_a;
                    alu_operand_b = op_b;
                end
            end
        end else begin
            always_comb begin
                op_a_sign_ext = op_a | ({AXI_ALU_RATIO*RISCV_WORD_WIDTH{sign_a}} & ~strb_ext);
                op_b_sign_ext = op_b | ({AXI_ALU_RATIO*RISCV_WORD_WIDTH{sign_b}} & ~strb_ext);

                if (atop_q[2:0] == axi_pkg::ATOP_SMAX || atop_q[2:0] == axi_pkg::ATOP_SMIN) begin
                    // Sign extend
                    alu_operand_a = op_a_sign_ext[addr_q[$clog2(AXI_DATA_WIDTH/8)-1:$clog2(RISCV_WORD_WIDTH/8)]];
                    alu_operand_b = op_b_sign_ext[addr_q[$clog2(AXI_DATA_WIDTH/8)-1:$clog2(RISCV_WORD_WIDTH/8)]];
                end else begin
                    // No sign extension necessary
                    alu_operand_a = op_a[addr_q[$clog2(AXI_DATA_WIDTH/8)-1:$clog2(RISCV_WORD_WIDTH/8)]];
                    alu_operand_b = op_b[addr_q[$clog2(AXI_DATA_WIDTH/8)-1:$clog2(RISCV_WORD_WIDTH/8)]];
                end
                res = '0;
                res[addr_q[$clog2(AXI_DATA_WIDTH/8)-1:$clog2(RISCV_WORD_WIDTH/8)]] = alu_result;
            end
        end
    endgenerate

    generate
        for (genvar i = 0; i < AXI_STRB_WIDTH; i++) begin
            always_comb begin
                if (strb_q[i]) begin
                    strb_ext[i] = 8'hFF;
                end else begin
                    strb_ext[i] = 8'h00;
                end
            end
        end
    endgenerate

    axi_riscv_amos_alu #(
        .DATA_WIDTH ( RISCV_WORD_WIDTH )
    ) i_amo_alu (
        .amo_op_i           ( atop_q        ),
        .amo_operand_a_i    ( alu_operand_a ),
        .amo_operand_b_i    ( alu_operand_b ),
        .amo_result_o       ( alu_result    )
    );

    // Validate parameters.
// pragma translate_off
`ifndef VERILATOR
    initial begin: validate_params
        assert (AXI_ADDR_WIDTH > 0)
            else $fatal(1, "AXI_ADDR_WIDTH must be greater than 0!");
        assert (AXI_DATA_WIDTH > 0)
            else $fatal(1, "AXI_DATA_WIDTH must be greater than 0!");
        assert (AXI_ID_WIDTH > 0)
            else $fatal(1, "AXI_ID_WIDTH must be greater than 0!");
        assert (AXI_MAX_WRITE_TXNS > 0)
            else $fatal(1, "AXI_MAX_WRITE_TXNS must be greater than 0!");
        assert (RISCV_WORD_WIDTH == 32 || RISCV_WORD_WIDTH == 64)
            else $fatal(1, "RISCV_WORD_WIDTH must be 32 or 64!");
        assert (RISCV_WORD_WIDTH <= AXI_DATA_WIDTH)
            else $fatal(1, "RISCV_WORD_WIDTH must not be greater than AXI_DATA_WIDTH!");
    end
`endif
// pragma translate_on

endmodule
